module top (
  input  logic  i,
  output logic  o 
);

assign o = i;

endmodule
